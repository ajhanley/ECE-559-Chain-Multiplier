module matrixReg(x, y, z);
//Matrix Register Holds x, horizontal dimension, y, the vertical dimension, and z, the actual matrixReg
	input[7:0] x,y;
	reg[x,y][7:0] matrix;//x by y 8 bit integers.




endmodule